(* SC_MODULE_EXPORT 	*)
module generator
(
 input clk,
 input enable,
 output [31:0] out
);
endmodule
